module ControlUnit();
    
endmodule