module EXE();

endmodule