module top()


endmodule