module MEM();



endmodule