module ID();


endmodule