module EXE();
    
endmodule