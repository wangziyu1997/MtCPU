module ID();
    ControlUnit cu ();
    regfile rf (inst[25:21],inst[20:16],res,wn,we,clock,resetn,ra,data);
    mux4 


endmodule