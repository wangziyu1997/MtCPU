module WB();
    
endmodule